//======================================================================
//  plate_cnn_fpga_top.v   –  all-in-one RTL for licence-plate CNN demo
//  • UART   : 115 200 baud, 8-N-1
//  • In     : 28×28  unsigned pixels  (784 bytes)
//
//  • Out    : 26×26  unsigned pixels  (676 bytes = first-layer feature map)
//              (pixel order: raster-scan)
//
//  Dependencies:
//     • weights.mem  (generated by export_weights.py)
//======================================================================

`timescale 1ns/1ps
//--------------------------------------------------------------------
//  Change these two parameters to match your board
//--------------------------------------------------------------------
`define CLK_HZ   12_000_000
`define BAUD     115200

//====================================================================
//  UART 8-N-1 Receiver  (unchanged from your uart_rx.sv)
//====================================================================
module uart_rx #(
    parameter CLK_HZ = `CLK_HZ,
    parameter BAUD   = `BAUD
)(
    input  wire clk,          // system clock
    input  wire rx,           // asynchronous serial in
    output reg  [7:0] data,   // received byte
    output reg        valid   // 1-clk pulse
);
    localparam DIV = CLK_HZ / BAUD;
    reg [$clog2(DIV)-1:0] cnt;
    reg [3:0] bitp;
    reg [7:0] sh;
    typedef enum logic [1:0] {IDLE,SRT,DATA,STP} state_t;
    state_t st /* synthesis syn_encoding = "onehot" */;

    always_ff @(posedge clk) begin
        valid <= 1'b0;
        case (st)
        IDLE: if (!rx) begin cnt <= DIV/2; st <= SRT; end
        SRT : if (!cnt--) begin cnt <= DIV-1; bitp <= 0; st <= DATA; end
        DATA: if (!cnt--) begin
                  cnt <= DIV-1;
                  sh  <= {rx, sh[7:1]};
                  if (bitp == 4'd7) st <= STP; else bitp <= bitp + 1'b1;
              end
        STP : if (!cnt--) begin data <= sh; valid <= 1'b1; st <= IDLE; end
        endcase
    end
endmodule

//====================================================================
//  UART 8-N-1 Transmitter  (unchanged from uart_tx.sv)
//====================================================================
module uart_tx #(
    parameter CLK_HZ = `CLK_HZ,
    parameter BAUD   = `BAUD
)(
    input  wire clk,
    input  wire [7:0] data,   // byte to send
    input  wire       valid,  // strobe 1 clk
    output wire       tx,     // serial data out
    output reg        busy    // 1 while shifting
);
    localparam DIV = CLK_HZ / BAUD;
    reg [$clog2(DIV)-1:0] cnt;
    reg [3:0] bitp;
    reg [9:0] sh;

    always_ff @(posedge clk) begin
        if (!busy && valid) begin
            sh   <= {1'b1, data, 1'b0};  // stop, data[7:0], start
            cnt  <= DIV-1;
            bitp <= 0;
            busy <= 1'b1;
        end else if (busy && !cnt--) begin
            cnt <= DIV-1;
            bitp <= bitp + 1'b1;
            if (bitp == 4'd9) busy <= 1'b0;
        end
        if (busy) sh <= {1'b1, sh[9:1]};
    end
    assign tx = busy ? sh[0] : 1'b1;
endmodule

//====================================================================
//  Weight ROM  (32 filters × 9 coeffs)     –  uses $readmemh
//====================================================================
module weight_rom #(parameter FILTS = 32)(
    input  wire [4:0] addr,                   // selects filter 0-31
    output reg  [8*9-1:0] data                // packed 9 × signed[7:0]
);
    reg [7:0] rom [0:FILTS-1][0:8];
    initial $readmemh("weights.mem", rom);

    always @* begin
        data = {
            rom[addr][0], rom[addr][1], rom[addr][2],
            rom[addr][3], rom[addr][4], rom[addr][5],
            rom[addr][6], rom[addr][7], rom[addr][8]
        };
    end
endmodule

//====================================================================
//  3×3 Sliding-window Conv2D   (verbatim from your conv2d_sliding.sv)
//  Note: this demo version stores the entire 5×5 image, suitable for
//        functional proof-of-concept. For production you would use a
//        line-buffer streaming core.
//====================================================================
module conv2d_sliding (
    input  wire clk,
    input  wire rst,
    input  wire start,
    input  wire [7:0] in_data,
    input  wire [7:0] kernel [0:8],   // 3×3 weights
    output reg  [15:0] out_data,
    output reg        done
);
    reg [7:0] input_buffer [0:24];  // 5×5 image (for demo)
    reg [5:0] in_idx;
    reg [3:0] out_idx;
    reg load_done, compute;

    integer sum;
    integer row, col, i, j;
    integer index;

    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            in_idx     <= 0;
            out_idx    <= 0;
            load_done  <= 0;
            compute    <= 0;
            done       <= 0;
        end else if (start && !load_done) begin
            input_buffer[in_idx] <= in_data;
            in_idx  <= in_idx + 1'b1;
            if (in_idx == 6'd24) begin
                load_done <= 1'b1;
                compute   <= 1'b1;
                out_idx   <= 0;
            end
        end else if (compute && out_idx < 9) begin
            row = out_idx / 3;
            col = out_idx % 3;
            sum = 0;
            for (i = 0; i < 3; i = i + 1) begin
                for (j = 0; j < 3; j = j + 1) begin
                    index = (row + i) * 5 + (col + j);
                    sum  += input_buffer[index] * kernel[i * 3 + j];
                end
            end
            out_data <= sum[15:0];
            out_idx  <= out_idx + 1'b1;
            if (out_idx == 3'd8)
                done <= 1'b1;
        end
    end
endmodule

//====================================================================
//  Top-level glue:  UART <--> Conv2D   (streaming 28×28 input)
//====================================================================
module plate_cnn_fpga_top (
    input  wire clk,
    input  wire rst_n,          // active-low
    input  wire uart_rx_i,
    output wire uart_tx_o
);
    //----------------------------------------------------------------
    //  (1) UART RX: receive 784 bytes – one 28×28 glyph
    //----------------------------------------------------------------
    wire [7:0] rx_byte;
    wire       rx_vld;
    uart_rx #(.CLK_HZ(`CLK_HZ), .BAUD(`BAUD)) RX (
        .clk(clk), .rx(uart_rx_i),
        .data(rx_byte), .valid(rx_vld)
    );

    //----------------------------------------------------------------
    //  (2) Weight ROM – we cycle through filter 0 only (demo)
    //----------------------------------------------------------------
    wire [8*9-1:0] kpacked;
    weight_rom ROM(.addr(5'd0), .data(kpacked));
    wire [7:0] kernel[0:8];
    genvar gi;
    generate
        for (gi=0; gi<9; gi=gi+1)
            assign kernel[gi] = kpacked[gi*8 +: 8];
    endgenerate

    //----------------------------------------------------------------
    //  (3) Simple state machine to feed conv2d_sliding demo core
    //----------------------------------------------------------------
    reg        start_d;
    reg [9:0]  byte_cnt;
    wire       conv_done;
    wire [15:0] conv_out;

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            byte_cnt <= 0;
            start_d  <= 0;
        end else if (rx_vld) begin
            byte_cnt <= byte_cnt + 1'b1;
            start_d  <= 1'b1;
        end else begin
            start_d  <= 1'b0;
        end
    end

    conv2d_sliding CONV (
        .clk   (clk),
        .rst   (~rst_n),
        .start (start_d),
        .in_data(rx_byte),
        .kernel(kernel),
        .out_data(conv_out),
        .done  (conv_done)
    );

    //----------------------------------------------------------------
    //  (4) UART TX: transmit the 9 conv results when done (demo)
    //----------------------------------------------------------------
    reg [7:0] tx_buf;
    reg       tx_req;
    reg [3:0] send_idx;

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            tx_req   <= 1'b0;
            send_idx <= 0;
        end else if (conv_done && send_idx < 9) begin
            tx_buf   <= conv_out[7:0];   // send LSB only for demo
            tx_req   <= 1'b1;
            send_idx <= send_idx + 1'b1;
        end else begin
            tx_req <= 1'b0;
        end
    end

    wire tx_busy;
    uart_tx #(.CLK_HZ(`CLK_HZ), .BAUD(`BAUD)) TX (
        .clk(clk), .data(tx_buf), .valid(tx_req),
        .busy(tx_busy), .tx(uart_tx_o)
    );

endmodule
